// Verilog module for Conway's Game of Life 16x16
