// Verilog module for Rule 90
