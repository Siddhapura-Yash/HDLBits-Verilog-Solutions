// Verilog module for Rule 110
